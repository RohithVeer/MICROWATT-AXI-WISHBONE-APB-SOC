/* Temporary stub: wb_to_apb.sv
   This file is a placeholder so the simulator can elaborate.
   Replace with the real implementation when available.
*/
module wb_to_apb (
  // generic ports — adjust or add ports if tests expect specific signals
  input  logic clk,
  input  logic rst_n
);
  // no behavior — stub only
endmodule
